.title nor_3_inp
.include techfile130.txt

vdd vdd 0 1.2

vA A 0 PULSE(0 1.2 2NS 2NS 2NS 50NS 100NS)
vB B 0 PULSE(0 1.2 20NS 2NS 2NS 50NS 100NS)
vC C 0 PULSE(0 1.2 30NS 2NS 2NS 50NS 100NS)

Mp1 1 A vdd vdd pmos l=120n w=8640n
Mp2 2 B 1 vdd pmos l=120n w=8640n
Mp3 vout C 2 vdd pmos l=120n w=8640n

Mn1 vout A 0 0 nmos l=120n w=960n
Mn2 vout B 0 0 nmos l=120n w=960n
Mn3 vout C 0 0 nmos l=120n w=960n


.tran 0.1n 200n 0 0.1n

.control
run 
plot v(A) v(B) v(vout)
.endc
.end
